module env

pub struct World {
mut:
	tiles [][]Tile
	cursor_x int
	curosr_y int
}