module main

fn main() {
	
}